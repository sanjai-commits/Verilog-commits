module helloWorld
  $display("Sanjai")
endmodule
